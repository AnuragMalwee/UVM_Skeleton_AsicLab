//Bock that encapsulates signals

interface our_interface(); 

    logic [7:0] input_1; //input_1
    logic [7:0] input_2; //input_2

    logic [15:0] output_3; //output

endinterface 